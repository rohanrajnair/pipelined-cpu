`include "mem.v"
`include "mux.v"
`include "alu.v"
`include "buff-1.v"
`include "cpu.v"

module top();

typedef enum { NOP=4'h0, MAX, UNUSED, STORE, ADD, INC, NEG, SUB, J, BRZ, JM, BRN, UNUSED1, UNUSED2, LOAD, SAVE_PC } opcode_t;

reg clk;
reg reset; 
int count;

always 
   #1 clk <= !clk;

initial begin
   clk = 0; 
   reset = 1;
   #50;
   init_imem();
   init_rf();
   init_dmem(); 
   reset = 0;
   #50;
   #50;
end 

always @ (posedge clk)
   begin
      if (reset)
         count = 0;
      else
         count += 1;

      if (count >= 2000) begin
          $display ("finished simulation");
          $finish;
      end
   end


function init_imem();
    [31:0] instr [255:0];
    int j = 0;

    for (int i=0; i < 256; i++) begin
        instr[i] = {LOAD, 6'h3, 6'h01, 6'h3f, 10'h0}; //load contents of mem pointed by register 1 into register 3
        instr[i] = {4'h0, 6'h1, 6'hf, 6'h0, 10'h0}; //NOP
    end
    //instr[4] = {LOAD, 6'h3, 6'h01, 6'h3f, 10'h0}; //load contents of mem pointed by register 1 into register 3
    //instr[4] = {SAVE_PC, 6'h3, 6'h01, 6'h3f, 10'h0}; //write 'h07f+pc(4) =='h83 into register 3
    //instr[4] = {STORE, 6'h6, 6'h05, 6'h4, 10'h0}; //store content of register 4 into [r5]
    //instr[24] = {INC, 6'h9, 6'h05, 6'h4, 10'h0}; //increment content of r5 into r9
    //instr[4] = {ADD, 6'h6, 6'h05, 6'h4, 10'h0}; //add register 4 & 5 into register 6
    //instr[32] = {BRZ, 6'h3, 6'h8, 6'h1, 10'h0}; //pc should NOT jump to 8
    //instr[36] = {NEG, 6'h6, 6'h05, 6'h4, 10'h0}; //twos complement of 5 into register 6
    //instr[40] = {SUB, 6'h6, 6'h07, 6'h4, 10'h0}; //r7-r4 into r6
    //instr[44] = {SUB, 6'h8, 6'h04, 6'h7, 10'h0}; //r4-r7 into r8. Should assert N at ALU as well
    //instr[48] = {SUB, 6'hA, 6'h04, 6'h4, 10'h0}; //r4-r4 into r10. Should assert Z at ALU as well
    //instr[48] = {J, 6'h3, 6'h2, 6'h1, 10'h0}; //pc should jump to 2
    //instr[52] = {BRZ, 6'h3, 6'h7, 6'h1, 10'h0}; //pc should jump to 7
    //instr[52] = {BRN, 6'h3, 6'h7, 6'h1, 10'h0}; //pc should NOT jump to 7
    //instr[56] = {SUB, 6'h8, 6'h04, 6'h7, 10'h0}; //r4-r7 into r8. Should assert N at ALU as well
    //instr[60] = {BRN, 6'h3, 6'h7, 6'h1, 10'h0}; //pc should jump to 7
    //instr[64] = {JM, 6'h3, 6'h2, 6'h1, 10'h0}; //pc should jump to 2
    

    //demo
   /*
    instr[j++] = {4'b1111, 6'b000001, 6'b000011, 6'b111111, 10'b0000000000}; //LDPC R1, 0xFF
    instr[j++] = {4'b0000, 6'b000000, 6'b000000, 6'b000000, 10'b0000000000}; //NOP
    instr[j++] = {4'b0000, 6'b000000, 6'b000000, 6'b000000, 10'b0000000000}; //NOP
    instr[j++] = {4'b0000, 6'b000000, 6'b000000, 6'b000000, 10'b0000000000}; //NOP
    instr[j++] = {4'b0101, 6'b000010, 6'b000001, 6'b000000, 10'b0000000000}; //INC R2, R1
    instr[j++] = {4'b0000, 6'b000000, 6'b000000, 6'b000000, 10'b0000000000}; //NOP
    instr[j++] = {4'b0000, 6'b000000, 6'b000000, 6'b000000, 10'b0000000000}; //NOP
    instr[j++] = {4'b0000, 6'b000000, 6'b000000, 6'b000000, 10'b0000000000}; //NOP

    instr[j++] = {4'b0110, 6'b000011, 6'b000001, 6'b000000, 10'b0000000000};  //NEG R3, R1
    instr[j++] = {4'b0000, 6'b000000, 6'b000000, 6'b000000, 10'b0000000000};  //NOP
    instr[j++] = {4'b0000, 6'b000000, 6'b000000, 6'b000000, 10'b0000000000}; //NOP
    instr[j++] = {4'b0000, 6'b000000, 6'b000000, 6'b000000, 10'b0000000000}; //NOP
    instr[j++] = {4'b1111, 6'b001010, 6'b000000, 6'b010010, 10'b0000000000}; //LDPC + 18
    instr[j++] = {4'b0000, 6'b000000, 6'b000000, 6'b000000, 10'b0000000000}; //NOP
    instr[j++] = {4'b0000, 6'b000000, 6'b000000, 6'b000000, 10'b0000000000}; //NOP
    instr[j++] = {4'b0000, 6'b000000, 6'b000000, 6'b000000, 10'b0000000000}; //NOP

    instr[j++] = {4'b1011, 6'b000000, 6'b001010, 6'b000000, 10'b0000000000}; //BRN R10
    instr[j++] = {4'b0000, 6'b000000, 6'b000000, 6'b000000, 10'b0000000000}; //NOP
    instr[j++] = {4'b0000, 6'b000000, 6'b000000, 6'b000000, 10'b0000000000}; //NOP
    instr[j++] = {4'b0000, 6'b000000, 6'b000000, 6'b000000, 10'b0000000000}; //NOP
    instr[j++] = {4'b0000, 6'b000000, 6'b000000, 6'b000000, 10'b0000000000}; //NOP
    instr[j++] = {4'b0101, 6'b000010, 6'b000010, 6'b000000, 10'b0000000000}; //INC R2, R2 (not taken)
    instr[j++] = {4'b0000, 6'b000000, 6'b000000, 6'b000000, 10'b0000000000}; //NOP
    instr[j++] = {4'b0000, 6'b000000, 6'b000000, 6'b000000, 10'b0000000000}; //NOP
    instr[j++] = {4'b0000, 6'b000000, 6'b000000, 6'b000000, 10'b0000000000}; //NOP


    //LABEL 1
    j = 30;

    instr[j++] = {4'b0011, 6'b000000, 6'b000001, 6'b000001, 10'b0000000000}; //ST R1, R1
    instr[j++] = {4'b0000, 6'b000000, 6'b000000, 6'b000000, 10'b0000000000}; //NOP
    instr[j++] = {4'b0000, 6'b000000, 6'b000000, 6'b000000, 10'b0000000000}; //NOP
    instr[j++] = {4'b0000, 6'b000000, 6'b000000, 6'b000000, 10'b0000000000}; //NOP
    instr[j++] = {4'b1110, 6'b000100, 6'b000001, 6'b000000, 10'b0000000000}; //LD R4, R1
    instr[j++] = {4'b0000, 6'b000000, 6'b000000, 6'b000000, 10'b0000000000}; //NOP
    instr[j++] = {4'b0000, 6'b000000, 6'b000000, 6'b000000, 10'b0000000000}; //NOP
    instr[j++] = {4'b0000, 6'b000000, 6'b000000, 6'b000000, 10'b0000000000}; //NOP
    instr[j++] = {4'b0100, 6'b000101, 6'b000001, 6'b000010, 10'b0000000000}; //ADD R5, R4, R1
    instr[j++] = {4'b0000, 6'b000000, 6'b000000, 6'b000000, 10'b0000000000}; //NOP
    instr[j++] = {4'b0000, 6'b000000, 6'b000000, 6'b000000, 10'b0000000000}; //NOP
    instr[j++] = {4'b0000, 6'b000000, 6'b000000, 6'b000000, 10'b0000000000}; //NOP
    instr[j++] = {4'b0111, 6'b000110, 6'b000100, 6'b000001, 10'b0000000000}; //SUB R6, R4, R1
    instr[j++] = {4'b0000, 6'b000000, 6'b000000, 6'b000000, 10'b0000000000}; //NOP
    instr[j++] = {4'b0000, 6'b000000, 6'b000000, 6'b000000, 10'b0000000000}; //NOP
    instr[j++] = {4'b0000, 6'b000000, 6'b000000, 6'b000000, 10'b0000000000}; //NOP
    instr[j++] = {4'b1111, 6'b001011, 6'b000000, 6'b001010, 10'b0000000000}; //LDPC + 14
    instr[j++] = {4'b0000, 6'b000000, 6'b000000, 6'b000000, 10'b0000000000}; //NOP
    instr[j++] = {4'b0000, 6'b000000, 6'b000000, 6'b000000, 10'b0000000000}; //NOP
    instr[j++] = {4'b0000, 6'b000000, 6'b000000, 6'b000000, 10'b0000000000}; //NOP
    instr[j++] = {4'b1001, 6'b000000, 6'b001011, 6'b000000, 10'b0000000000}; //BRZ R11
    instr[j++] = {4'b0000, 6'b000000, 6'b000000, 6'b000000, 10'b0000000000}; //NOP
    instr[j++] = {4'b0000, 6'b000000, 6'b000000, 6'b000000, 10'b0000000000}; //NOP
    instr[j++] = {4'b0000, 6'b000000, 6'b000000, 6'b000000, 10'b0000000000}; //NOP
    instr[j++] = {4'b0000, 6'b000000, 6'b000000, 6'b000000, 10'b0000000000}; //NOP
    instr[j++] = {4'b0101, 6'b000010, 6'b000010, 6'b000000, 10'b0000000000}; //INC R2, R2
    instr[j++] = {4'b0000, 6'b000000, 6'b000000, 6'b000000, 10'b0000000000}; //NOP
    instr[j++] = {4'b0000, 6'b000000, 6'b000000, 6'b000000, 10'b0000000000}; //NOP
    instr[j++] = {4'b0000, 6'b000000, 6'b000000, 6'b000000, 10'b0000000000}; //NOP

    j = 60;
    //LABEL 2
    instr[60] = {4'b1010, 6'b000000, 6'b000001, 6'b000000, 10'b0000000000}; //JM R1
    instr[61] = {4'b0000, 6'b000000, 6'b000000, 6'b000000, 10'b0000000000}; //NOP
    instr[62] = {4'b0000, 6'b000000, 6'b000000, 6'b000000, 10'b0000000000}; //NOP
    instr[63] = {4'b0000, 6'b000000, 6'b000000, 6'b000000, 10'b0000000000}; //NOP


    j = 255;
   //OXFF:
   instr[255] = {4'b1000, 6'b000000, 6'b000001, 6'b000000, 10'b0000000000}; //J R1
   instr[256] = {4'b0000, 6'b000000, 6'b000000, 6'b000000, 10'b0000000000}; //NOP
   instr[257] = {4'b0000, 6'b000000, 6'b000000, 6'b000000, 10'b0000000000}; //NOP
   instr[258] = {4'b0000, 6'b000000, 6'b000000, 6'b000000, 10'b0000000000}; //NOP
   */
  
  
  //max function  
  
   instr[0] = {4'b1110, 6'b000000, 6'b000001, 6'b000000, 10'b0000000000}; // LOAD R0, R1
   instr[1] = {4'b0000, 6'b000000, 6'b000000, 6'b000000, 10'b0000000000}; // NOP
   instr[2] = {4'b0000, 6'b000000, 6'b000000, 6'b000000, 10'b0000000000}; // NOP
   instr[3] = {4'b0000, 6'b000000, 6'b000000, 6'b000000, 10'b0000000000}; // NOP
   instr[4] = {4'b0000, 6'b000000, 6'b000000, 6'b000000, 10'b0000000000}; // NOP
   instr[5] = {4'b1000, 6'b000000, 6'b010100, 6'b000000, 10'b0000000000}; // J LOOP
   instr[6] = {4'b0000, 6'b000000, 6'b000000, 6'b000000, 10'b0000000000}; // NOP
   instr[7] = {4'b0000, 6'b000000, 6'b000000, 6'b000000, 10'b0000000000}; // NOP
   instr[8] = {4'b0000, 6'b000000, 6'b000000, 6'b000000, 10'b0000000000}; // NOP
   instr[9] = {4'b0000, 6'b000000, 6'b000000, 6'b000000, 10'b0000000000}; // NOP
   
   // LOOP
   instr[20] = {4'b1001, 6'b000000, 6'b010101, 6'b000000, 10'b0000000000}; // BRZ END
   instr[21] = {4'b0000, 6'b000000, 6'b000000, 6'b000000, 10'b0000000000}; // NOP
   instr[22] = {4'b0000, 6'b000000, 6'b000000, 6'b000000, 10'b0000000000}; // NOP
   instr[23] = {4'b0000, 6'b000000, 6'b000000, 6'b000000, 10'b0000000000}; // NOP
   instr[24] = {4'b0000, 6'b000000, 6'b000000, 6'b000000, 10'b0000000000}; // NOP
   instr[25] = {4'b0100, 6'b000001, 6'b000001, 6'b011110, 10'b0000000000}; // ADD R1, R1, R30
   instr[26] = {4'b0000, 6'b000000, 6'b000000, 6'b000000, 10'b0000000000}; // NOP
   instr[27] = {4'b0000, 6'b000000, 6'b000000, 6'b000000, 10'b0000000000}; // NOP
   instr[28] = {4'b0000, 6'b000000, 6'b000000, 6'b000000, 10'b0000000000}; // NOP
   instr[29] = {4'b0000, 6'b000000, 6'b000000, 6'b000000, 10'b0000000000}; // NOP
   instr[30] = {4'b1110, 6'b000111, 6'b000001, 6'b000000, 10'b0000000000}; //LOAD R7, R1
   instr[31] = {4'b0000, 6'b000000, 6'b000000, 6'b000000, 10'b0000000000}; // NOP
   instr[32] = {4'b0000, 6'b000000, 6'b000000, 6'b000000, 10'b0000000000}; // NOP
   instr[33] = {4'b0000, 6'b000000, 6'b000000, 6'b000000, 10'b0000000000}; // NOP
   instr[34] = {4'b0000, 6'b000000, 6'b000000, 6'b000000, 10'b0000000000}; // NOP
   
   
   
   instr[35] = {4'b0111, 6'b001001, 6'b000000, 6'b000111, 10'b0000000000}; // SUB R9, R0, R7
   instr[36] = {4'b0000, 6'b000000, 6'b000000, 6'b000000, 10'b0000000000}; // NOP
   instr[37] = {4'b0000, 6'b000000, 6'b000000, 6'b000000, 10'b0000000000}; // NOP
   instr[38] = {4'b0000, 6'b000000, 6'b000000, 6'b000000, 10'b0000000000}; // NOP
   instr[39] = {4'b0000, 6'b000000, 6'b000000, 6'b000000, 10'b0000000000}; // NOP
   instr[40] = {4'b1011, 6'b000000, 6'b010110, 6'b000000, 10'b0000000000}; // BRN IF
   instr[41] = {4'b0000, 6'b000000, 6'b000000, 6'b000000, 10'b0000000000}; // NOP
   instr[42] = {4'b0000, 6'b000000, 6'b000000, 6'b000000, 10'b0000000000}; // NOP
   instr[43] = {4'b0000, 6'b000000, 6'b000000, 6'b000000, 10'b0000000000}; // NOP
   instr[44] = {4'b0000, 6'b000000, 6'b000000, 6'b000000, 10'b0000000000}; // NOP
   instr[45] = {4'b0111, 6'b000010, 6'b000010, 6'b011110, 10'b0000000000}; // SUB R2, R2, R30
   instr[46] = {4'b0000, 6'b000000, 6'b000000, 6'b000000, 10'b0000000000}; // NOP
   instr[47] = {4'b0000, 6'b000000, 6'b000000, 6'b000000, 10'b0000000000}; // NOP
   instr[48] = {4'b0000, 6'b000000, 6'b000000, 6'b000000, 10'b0000000000}; // NOP
   instr[49] = {4'b0000, 6'b000000, 6'b000000, 6'b000000, 10'b0000000000}; // NOP
   instr[50] = {4'b1000, 6'b000000, 6'b010100, 6'b000000, 10'b0000000000}; // J LOOP
   instr[51] = {4'b0000, 6'b000000, 6'b000000, 6'b000000, 10'b0000000000}; // NOP
   instr[52] = {4'b0000, 6'b000000, 6'b000000, 6'b000000, 10'b0000000000}; // NOP
   instr[53] = {4'b0000, 6'b000000, 6'b000000, 6'b000000, 10'b0000000000}; // NOP
   instr[54] = {4'b0000, 6'b000000, 6'b000000, 6'b000000, 10'b0000000000}; // NOP
   
   // IF
   
   instr[60] = {4'b0100, 6'b000000, 6'b000111, 6'b011111, 10'b0000000000}; // ADD R0, R7, R31
   instr[61] = {4'b0000, 6'b000000, 6'b000000, 6'b000000, 10'b0000000000}; // NOP
   instr[62] = {4'b0000, 6'b000000, 6'b000000, 6'b000000, 10'b0000000000}; // NOP
   instr[63] = {4'b0000, 6'b000000, 6'b000000, 6'b000000, 10'b0000000000}; // NOP
   instr[64] = {4'b0000, 6'b000000, 6'b000000, 6'b000000, 10'b0000000000}; // NOP
   instr[65] = {4'b0111, 6'b000010, 6'b000010, 6'b011110, 10'b0000000000}; // SUB R2, R2, R30
   instr[66] = {4'b0000, 6'b000000, 6'b000000, 6'b000000, 10'b0000000000}; // NOP
   instr[67] = {4'b0000, 6'b000000, 6'b000000, 6'b000000, 10'b0000000000}; // NOP
   instr[68] = {4'b0000, 6'b000000, 6'b000000, 6'b000000, 10'b0000000000}; // NOP
   instr[69] = {4'b0000, 6'b000000, 6'b000000, 6'b000000, 10'b0000000000}; // NOP
   instr[70] = {4'b1000, 6'b000000, 6'b010100, 6'b000000, 10'b0000000000}; // J LOOP
   instr[71] = {4'b0000, 6'b000000, 6'b000000, 6'b000000, 10'b0000000000}; // NOP
   instr[72] = {4'b0000, 6'b000000, 6'b000000, 6'b000000, 10'b0000000000}; // NOP
   instr[73] = {4'b0000, 6'b000000, 6'b000000, 6'b000000, 10'b0000000000}; // NOP
   instr[74] = {4'b0000, 6'b000000, 6'b000000, 6'b000000, 10'b0000000000}; // NOP
      
  
  //max instruction
  // instr[0] = {4'b0001, 6'b000001, 6'b001010, 6'b001011, 10'b0000000000}; // MAX R1, R10, R11


    for (int i=0; i < 256; i++) begin
      cpu_inst.imem_inst.mem[i] = instr[i];
    end
endfunction

function init_rf();
   [31:0] register [63:0];

   for (bit[7:0] i =0; i < 8'd64; i++) begin
     register[i] = {i,i,i,i};
   end

   //max function
    
   register[0] = 32'd0;    
   register[1] = 32'd10;   // base address of A
   register[2] = 32'd6;    // # elements in A
   register[3] = 32'b1;    // i 
   register[20] = 32'd20;  // loop label
   register[21] = 32'd50;  // end label
   register[22] = 32'd60;  // if label
   register[30] = 32'b1;
   register[31] = 32'b0;
   
   
   //max instruction
   //register[10] = 32'd50;
   //register[11] = 32'd4; 

   for (int i = 0; i < 64; i++) begin
      cpu_inst.rf_inst.mem[i] = register[i];
   end
endfunction


function init_dmem();
   [31:0] data [63:0];

   data[0] = 32'hb2301_0010;
   data[1] = 32'hb2101_0123;
   data[2] = 32'h0011_bae2;
   data[3] = 32'h0023_124b;

   data[10] = 32'd30; //A
   data[11] = 32'd8;
   data[12] = 32'd11;
   data[13] = 32'd18;
   data[14] = 32'd 60;
   data[15] = 32'd 40; 

   //max instruction
   data[50] = 32'd45;
   data[51] = 32'd20;
   data[52] = 32'd70;
   data[53] = 32'd5;


   for (int i = 0; i < 2**16; i++) begin
      cpu_inst.dmem_inst.mem[i] = data[i];
   end


endfunction



cpu cpu_inst(.clk(clk),
             .reset(reset)
);


endmodule 
